library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
entity dsp_1 is
Port ( clk : in STD_LOGIC;
sin : in STD_LOGIC;
din : in STD_LOGIC_VECTOR (23 downto 0);
dout : out STD_LOGIC_VECTOR (23 downto 0));
end dsp_1;
architecture Behavioral of dsp_1 is
component koefmem is port(
clka : IN std_logic;
addra : IN std_logic_vector(15 downto 0);
douta : OUT std_logic_vector(11 downto 0));
end component;
type firkoefmem is array(255 downto 0) of signed(17 downto 0);
signal dfir : firkoefmem := (
"100000000000000000", "011101010110001100", "010101111101111100", "001011011101001001", "000000000000000000", "110101110101111100",
"101110101111100101", "101011100111001010", "101100011001000000", "110000001100101000", "110101101010000010", "111011010100001010",
"000000000000000000", "000011000011000101", "000100010110010010", "000100001110101101", "000011010000101000", "000010000001011100",
"000000111101001101", "000000010001110100", "000000000000000000", "111111111111111011", "000000000111001010", "000000001101011100",
"000000001110110101", "000000001011100100", "000000000110010100", "000000000001111010", "000000000000000000", "000000000000011111",
"000000000010001100", "000000000011101001", "000000000011111110", "000000000011000111", "000000000001101100", "000000000000011110",
"000000000000000000", "000000000000010000", "000000000000111001", "000000000001011011", "000000000001100010", "000000000001001101",
"000000000000101001", "000000000000001010", "000000000000000000", "000000000000001001", "000000000000011100", "000000000000101100",
"000000000000101111", "000000000000100100", "000000000000010011", "000000000000000100", "000000000000000000", "000000000000000101",
"000000000000001111", "000000000000011000", "000000000000011001", "000000000000010011", "000000000000001010", "000000000000000010",
"000000000000000000", "000000000000000011", "000000000000001001", "000000000000001110", "000000000000001111", "000000000000001011",
"000000000000000110", "000000000000000001", "000000000000000000", "000000000000000010", "000000000000000110", "000000000000001001",
"000000000000001001", "000000000000000111", "000000000000000011", "000000000000000000", "000000000000000000", "000000000000000001",
"000000000000000100", "000000000000000110", "000000000000000110", "000000000000000101", "000000000000000010", "000000000000000000",
"000000000000000000", "000000000000000001", "000000000000000011", "000000000000000100", "000000000000000100", "000000000000000011",
"000000000000000001", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000010", "000000000000000011",
"000000000000000011", "000000000000000010", "000000000000000001", "000000000000000000", "000000000000000000", "000000000000000000",
"000000000000000001", "000000000000000010", "000000000000000010", "000000000000000010", "000000000000000001", "000000000000000000",
"000000000000000000", "000000000000000000", "000000000000000001", "000000000000000001", "000000000000000010", "000000000000000001",
"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000001",
"000000000000000001", "000000000000000001", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
"000000000000000000", "000000000000000001", "000000000000000001", "000000000000000001", "000000000000000000", "000000000000000000",
"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000001", "000000000000000000",
"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000",
"000000000000000000", "000000000000000000", "000000000000000000", "000000000000000000");
type inputbank is array(255 downto 0) of signed(23 downto 0);
signal inputs : inputbank;
signal dct1 : signed(35 downto 0) := (others => '0');
signal dct2 : signed(36 downto 0) := (others => '0');
type dctbank is array(255 downto 0) of signed(26 downto 0);
signal dcts : dctbank;
signal fir1 : signed(44 downto 0) := (others => '0');
type firbank is array(255 downto 0) of signed(28 downto 0);
signal firs : firbank;
signal idct0 : signed(40 downto 0) := (others => '0');
signal idct1 : signed(40 downto 0) := (others => '0');
signal idct2 : signed(40 downto 0) := (others => '0');
signal idct3 : signed(23 downto 0) := (others => '0');
type idctbank is array(255 downto 0) of signed(23 downto 0);
signal idcts : idctbank:= (others => (others => '0'));
signal koef : std_logic_vector(11 downto 0) := (others => '0');
signal add : std_logic_vector(15 downto 0) := (others => '0');
signal addr : signed(16 downto 0):= (others => '0');
signal i, j, k, l : integer := 0;
signal en : std_logic := '0';
type statelist is (idle, io, dct, fir, idct, jeda);
signal state : statelist := idle;
begin
Koefisien:koefmem port map(clka => clk, addra => add, douta => koef);
Proses:process(clk, en, j, k, din, en, sin, dfir, koef)
begin
if rising_edge(clk) then
case state iswhen idle => if sin = '1' then
state <= io;
dout <= "000000000000000000000000";
end if;
when io =>if en = '1' then
if j < 257 then
if j = 256 then
state <= dct;
j <= 0;
else
inputs(j) <= signed(din);
dout <= std_logic_vector(idcts(j));
j <= j + 1;
end if;
end if;
end if;
when dct =>if j < 257 then
if j = 256 then
j <= 0;
addr <= (others => '0');
state <= fir;
else
if k < 257 then
if k = 256 then
k <= 0;
j <= j + 1;
dct2(36 downto 1) <= dct1;
dcts(j) <= dct2(36 downto 10);
elsif k = 0 then
addr <= addr + "00000000000000001";
dct1 <= signed(koef) * inputs(k);
k <= k + 1;
else
addr <= addr + "00000000000000001";
dct1 <= dct1 + signed(koef) * inputs(k);
k <= k + 1;
end if;
end if;
end if;
end if;
when fir =>
if k < 257 then
if k = 256 then
k <= 0;
j <= j + 1;
state <= idct;
elsif k = 0 then
fir1 <= dfir(k) * dcts(k);
firs(k) <= fir1(44 downto 16);
idct0 <= fir1(44 downto 4);
k <= k + 1;
else
fir1 <= dfir(k) * dcts(k);
firs(k) <= fir1(44 downto 16);
k <= k + 1;
end if;
end if;
when idct =>if j < 257 then
if j = 256 then
j <= 0;
addr <= (others => '0');
state <= jeda;
else
if k < 257 then
if k = 256 then
k <= 0;
j <= j + 1;
idct2 <= idct0 + idct1;
idct3(22 downto 0) <= idct2(40 downto 18);
idct3(23) <= idct2(40);
idcts(j) <= idct3;
elsif k = 0 then
addr <= addr + "00000000000000001";
idct1 <= signed(koef) * firs(k);
k <= k + 1;
else
addr <= addr + "00000000000000001";
idct1 <= idct1 + signed(koef) * firs(k);
k <= k + 1;
end if;
end if;
end if;
end if;
when jeda =>
if k < 124673 then
if k = 124673 then
k <= 0;
state <= idle;
else
k <= k + 1;
end if;
end if;
when others => state <= idle;
end case;
end if;
end process;
add <= std_logic_vector(addr(15 downto 0));
Enable:process(clk, i)
begin
if rising_edge(clk) then
if i < 1001 then
if i = 1000 then
i <= 0;
else
i <= i + 1;
en <= '0';
if i = 0 then
en <= '1';
end if;
end if;
end if;
end if;
end process;
end Behavioral;
